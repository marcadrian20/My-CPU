library verilog;
use verilog.vl_types.all;
entity BOARD_tb is
end BOARD_tb;
